interface intff;
  logic a, b, c;
  logic sum, carry;
endinterface
