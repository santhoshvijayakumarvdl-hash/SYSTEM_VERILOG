
class name;
  int a;
  bit b;
  
  function new ();
    a=5;
     b=1;
  endfunction
  
  
  
  function void display1();
    $display("%b %b ",a,b);
  endfunction
endclass


class name2 extends name;
  int c;
  bit d;
 
  
  function new();
    c=6;
     d=0;
 
  endfunction
  
  
  
  function void display();
    $display("%b %b %b %b",a,b,c,d);
  endfunction
endclass


module tb;
  initial begin
    name2 g1;
    g1=new();
    g1.display();
    g1.display1();
     
    

  end
endmodule
    
