interface intff;
  logic clk,rst;
  logic d,d_out;
endinterface
